* SPICE3 file created from inv_layout.ext - technology: sample_6m

.option scale=0.09u

M1000 out in vdd vdd cmosp w=8 l=2
+  ad=48 pd=28 as=48 ps=28
M1001 out in gnd gnd cmosn w=4 l=2
+  ad=29 pd=22 as=29 ps=22
